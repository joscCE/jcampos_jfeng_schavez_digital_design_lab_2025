module tb_TopDecoder();
	

endmodule